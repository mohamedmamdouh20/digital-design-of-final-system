
/////////////////////////////////////////////////////////////
/////////////////////// buffer			 ////////////////////////
/////////////////////////////////////////////////////////////

module buffer (
input      IN,
output     OUT
);

//buf buffer(OUT,IN);
CLKBUFX6M delay(.A(IN),.Y(OUT));



endmodule
